library verilog;
use verilog.vl_types.all;
entity computer_sim is
end computer_sim;
