library verilog;
use verilog.vl_types.all;
entity clock_sim is
end clock_sim;
